`timescale 1ns/1ps

/////////////
//
/////////////

module hilbert_control (
				input clock,
				input reset,
				input start,   // set to 1 for one clock to start 
				output enable,
				output reg [5:0] count

);

endmodule

